
module Sequential_TB();

//ToDo

endmodule